`timescale 1ns/1ns

module thermo_to_onehot(
    thermo,
    onehot
    );

// TO DO

endmodule
