`timescale 1ns/1ns

module onehot_to_bin(
    onehot,
    bin
    );

// TO DO

endmodule
