`timescale 1ns/1ns

module majority(
    in1,
    in2,
    in3,
    in4,
    out
    );

// TO DO

endmodule
