`timescale 1ns/1ns

module thermo_to_bin(
    thermo,
    bin
    );

// TO DO

endmodule
