`timescale 1ns/1ns

module tb_thermo_maj;

// TO DO

endmodule


