// Code your testbench here
// or browse Examples
`include "tb_thermo_maj.v"


